module top_dummy();
    initial begin
        $display("Project Initialized - Work In Progress");
        #10 $finish;
    end
endmodule
